// Test file for Verilog completion
module test_module(
    input wire clk,
    output reg data_out
);

// Type 'mod' and press Ctrl+Space to test completion
// Type 'al' and press Ctrl+Space to test completion
// Type 'reg' and press Ctrl+Space to test completion

endmodule